
//`include "checker.sv"
//`include "simple.sv"
//`include "soft_cstr.sv"
//`include "post_rand.sv"
//`include "post_count_ones.sv"
//`include "cstr_inheritance_polymorphis.sv"
//`include "cstr_inheritance_polymorphism_ex2.sv"
//`include "cstr_inheritance_ex1.sv"

