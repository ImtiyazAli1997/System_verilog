module tb;
	
	initial begin
	
		$display("Newyork is awesom place.
		So energitic and  vibrant");
	end
	
endmodule